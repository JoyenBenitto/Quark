// This is th etop module 

package quark;

    import regfile :: *;

    module mkquark;

    endmodule: mkquark

endpackage!