package Fn_Decode

import Instr_Bits :: * ;
import Inter_Stage :: * ;

endpackage: Fn_Decode