package Arch



endpackage
